      12          0.73707654          0.00034632  0.34576000          80    41.0   99   96.16
      16          1.23653117          0.00057169  0.34576000          80    41.0   99   97.87
      24          2.58120956          0.00117779  0.34576000          80    41.0   99   70.10
      32          4.36655847          0.00196474  0.34576000          80    41.0   99   94.39
      48          9.18873404          0.00407377  0.34576000          80    41.0   99  117.43
      64         15.64108214          0.00687892  0.34576000          80    41.0   99  106.39
      96         33.21421640          0.01427422  0.34576000          80    41.0   99   92.78
     128         56.86188056          0.02405585  0.34576000          80    41.0   99  111.49
     156         82.36380467          0.03467201  0.34576000          80    41.0   99  108.00
     198        128.99824202          0.05351899  0.34576000          80    41.0   99  103.01
     256        209.42477800          0.08522265  0.34576000          80    41.0   99   87.96
     512        785.85035377          4.17267171  0.34565000          80     0.2    0    0.00
